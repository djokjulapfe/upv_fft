library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity upv_fft is
	port (
		uart_in  : in  std_logic;
		uart_out : out std_logic
	);
end entity upv_fft;

architecture behav of upv_fft is
begin
end architecture behav;